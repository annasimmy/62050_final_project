module video_sig_gen
#(
  parameter ACTIVE_H_PIXELS = 1280,
  parameter H_FRONT_PORCH = 110,
  parameter H_SYNC_WIDTH = 40,
  parameter H_BACK_PORCH = 220,
  parameter ACTIVE_LINES = 720,
  parameter V_FRONT_PORCH = 5,
  parameter V_SYNC_WIDTH = 5,
  parameter V_BACK_PORCH = 20,
  parameter FPS = 60)
(
  input wire pixel_clk_in,
  input wire rst_in,
  output logic [$clog2(TOTAL_PIXELS)-1:0] hcount_out,
  output logic [$clog2(TOTAL_LINES)-1:0] vcount_out,
  output logic vs_out, //vertical sync out
  output logic hs_out, //horizontal sync out
  output logic ad_out, // active drawing
  output logic nf_out, //single cycle enable signal
  output logic [5:0] fc_out); //frame

  localparam TOTAL_LINES = ACTIVE_LINES + V_FRONT_PORCH + V_SYNC_WIDTH + V_BACK_PORCH; //figure this out
  localparam TOTAL_WIDTH = ACTIVE_H_PIXELS + H_FRONT_PORCH + H_SYNC_WIDTH + H_BACK_PORCH;
  localparam TOTAL_PIXELS = TOTAL_LINES * TOTAL_WIDTH; //figure this out

  
  //your code here
  always_ff @(posedge pixel_clk_in) begin
    if(rst_in) begin
      hcount_out <= 0;
      vcount_out <= 0;
      vs_out <= 0;
      hs_out <= 0;
      ad_out <= 0;
      nf_out <= 0;
      fc_out <= 0;
    end else begin
      if(hcount_out == 0 && vcount_out == 0 && !ad_out) begin
        ad_out <= 1;
      end else if(hcount_out + 1 == TOTAL_WIDTH) begin
        hcount_out <= 0;
        if(vcount_out + 1 == TOTAL_LINES) begin
          vcount_out <= 0;
          ad_out <= 1;
        end else begin
          vcount_out <= vcount_out + 1;
          hs_out <= 0;
          if(vcount_out + 1 >= ACTIVE_LINES + V_FRONT_PORCH && vcount_out + 1 < ACTIVE_LINES + V_FRONT_PORCH + V_SYNC_WIDTH) begin
            vs_out <= 1;
          end else begin
            vs_out <= 0;
            hs_out <= 0;
            ad_out <= 0;
          end
          if(vcount_out + 1 < ACTIVE_LINES) begin
            ad_out <= 1;
          end else begin
            ad_out <= 0;
          end
        end
      end else begin
        hcount_out <= hcount_out + 1;
        if(hcount_out + 1 >= ACTIVE_H_PIXELS + H_FRONT_PORCH && hcount_out + 1 < ACTIVE_H_PIXELS + H_FRONT_PORCH + H_SYNC_WIDTH) begin
          hs_out <= 1;
        end else begin
          hs_out <= 0;
        end
        if(vcount_out < ACTIVE_LINES && hcount_out + 1 < ACTIVE_H_PIXELS) begin
          ad_out <= 1;
        end else begin
          ad_out <= 0;
        end
        if(vcount_out == ACTIVE_LINES && hcount_out + 1 == ACTIVE_H_PIXELS) begin
          nf_out <= 1;
          if(fc_out == 59) begin
            fc_out <= 0;
          end else begin
            fc_out <= fc_out + 1;
          end
        end else begin
          nf_out <= 0;
        end
      end
    end
  end

endmodule